* Extracted by KLayout with GF180MCU LVS runset on : 15/02/2026 00:48

.SUBCKT NAND2 vdd OUT vss IN1 IN0
M$1 OUT IN1 vdd vdd pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$2 OUT IN0 vdd vdd pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$3 \$6 IN1 OUT vss nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$4 \$6 IN0 vss vss nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
.ENDS NAND2
