* NGSPICE file created from dff_flat.ext - technology: gf180mcuD

.subckt dff_flat RSTN VDD CLK VSS D Q Qb
X0 a_n249_n4912# a_n1374_n6642# a_991_n4911# VSS.t1 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X1 VSS.t13 a_n359_n5759.t3 Q.t0 VSS.t12 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X2 a_n359_n5759.t1 a_n249_n4912# VDD.t17 VDD.t16 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X3 VDD.t15 RSTN.t0 a_881_n5758# VDD.t14 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X4 VDD.t3 a_n1374_n6642# a_1067_n6116# VDD.t2 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X5 a_2281_n4424# D.t0 a_1056_n4015# VSS.t11 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X6 VSS.t10 CLK.t0 a_n1342_n5730# VSS.t9 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X7 a_2280_n3998# D.t1 a_1056_n4015# VDD.t13 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X8 VDD.t19 CLK.t1 a_n1342_n5730# VDD.t18 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X9 VSS.t24 a_n1342_n5730# a_n1374_n6642# VSS.t23 nfet_03v3 ad=0.2667p pd=2.11u as=0.2625p ps=2.09u w=0.42u l=0.28u
X10 a_1059_n5756# a_991_n4911# a_881_n5758# VSS.t25 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X11 VSS.t5 a_1056_n4015# a_991_n4911# VSS.t4 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X12 VSS.t22 a_n1342_n5730# a_1068_n6542# VSS.t21 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X13 VSS.t8 a_n912_n3722# Qb.t0 VSS.t7 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X14 VSS.t3 RSTN.t1 a_n181_n5757# VSS.t2 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X15 VDD.t12 a_n359_n5759.t4 Q.t1 VDD.t11 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X16 a_n249_n4912# a_n1342_n5730# a_991_n4911# VDD.t23 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X17 VSS.t16 a_n359_n5759.t5 a_n912_n3722# VSS.t15 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X18 VDD.t22 a_n1342_n5730# a_n1374_n6642# VDD.t21 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X19 a_881_n5758# a_n1374_n6642# a_1056_n4015# VSS.t0 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X20 VDD.t7 a_n912_n3722# Qb.t1 VDD.t6 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X21 VSS.t20 a_n1342_n5730# a_2281_n4424# VSS.t19 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X22 VDD.t27 RSTN.t2 a_n359_n5759.t2 VDD.t26 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X23 VDD.t1 a_n1374_n6642# a_2280_n3998# VDD.t0 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X24 a_1067_n6116# a_n359_n5759.t6 a_n249_n4912# VDD.t10 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X25 a_881_n5758# a_991_n4911# VDD.t25 VDD.t24 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X26 VSS.t18 RSTN.t3 a_1059_n5756# VSS.t17 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X27 VDD.t5 a_1056_n4015# a_991_n4911# VDD.t4 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X28 a_881_n5758# a_n1342_n5730# a_1056_n4015# VDD.t20 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X29 a_1068_n6542# a_n359_n5759.t7 a_n249_n4912# VSS.t6 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X30 a_n181_n5757# a_n249_n4912# a_n359_n5759.t0 VSS.t14 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X31 VDD.t9 a_n359_n5759.t8 a_n912_n3722# VDD.t8 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
R0 VSS.n23 VSS.n16 749278
R1 VSS.n16 VSS.t11 91327.6
R2 VSS.n5 VSS.n3 64653.5
R3 VSS.n50 VSS.n3 47027.8
R4 VSS.n13 VSS.n8 11150.5
R5 VSS.t7 VSS.n46 10656.3
R6 VSS.n46 VSS.n45 9310.54
R7 VSS.n6 VSS.n3 9172.39
R8 VSS.n17 VSS.n8 8859.18
R9 VSS.n46 VSS.n7 7710.44
R10 VSS.n43 VSS.n9 6769.51
R11 VSS.n35 VSS.n34 6625.47
R12 VSS.n45 VSS.n8 5874.35
R13 VSS.t23 VSS.n49 4464.13
R14 VSS.n13 VSS.n11 4354.26
R15 VSS.n30 VSS.n10 4226.8
R16 VSS.n29 VSS.n11 4102.23
R17 VSS.n45 VSS.n44 3676.98
R18 VSS.n24 VSS.n23 3564.92
R19 VSS.n44 VSS.t0 2894.81
R20 VSS.n47 VSS.n7 2588.74
R21 VSS.t12 VSS.n3 2474.65
R22 VSS.n49 VSS.n48 2224.45
R23 VSS.n49 VSS.t9 1774.36
R24 VSS.n48 VSS.n6 1755.92
R25 VSS.n22 VSS.n21 1702.15
R26 VSS.t4 VSS.n24 1689.9
R27 VSS.n24 VSS.n10 1589.78
R28 VSS.t9 VSS.n5 1493.57
R29 VSS.t19 VSS.n15 1430.46
R30 VSS.n25 VSS.t4 1413.04
R31 VSS.t25 VSS.n9 1360.03
R32 VSS.n21 VSS.t0 1205.49
R33 VSS.t15 VSS.n7 1196.19
R34 VSS.n48 VSS.n47 1177.13
R35 VSS.n18 VSS.t17 1172.44
R36 VSS.n23 VSS.n22 1095.11
R37 VSS.n25 VSS.n11 1090.87
R38 VSS.n36 VSS.t2 1070.49
R39 VSS.n34 VSS.t6 1055.67
R40 VSS.n42 VSS.t15 992.063
R41 VSS.n30 VSS.t1 940.115
R42 VSS.n50 VSS.t23 920.712
R43 VSS.t11 VSS.t19 915.494
R44 VSS.n18 VSS.n10 900.433
R45 VSS.n34 VSS.n33 836.077
R46 VSS.n36 VSS.n35 822.135
R47 VSS.n32 VSS.n30 797.649
R48 VSS.t17 VSS.t25 750.361
R49 VSS.t2 VSS.t14 685.112
R50 VSS.n17 VSS.n16 674.74
R51 VSS.n38 VSS.n7 671.655
R52 VSS.n43 VSS.n42 615.08
R53 VSS.n33 VSS.t12 604.99
R54 VSS.t21 VSS.n32 576.241
R55 VSS.t1 VSS.n29 492.724
R56 VSS.n44 VSS.n43 472.2
R57 VSS.n15 VSS.n13 469.19
R58 VSS.t14 VSS.n6 466.733
R59 VSS.n47 VSS.t7 415.238
R60 VSS.t6 VSS.t21 368.795
R61 VSS.n35 VSS.n9 317.529
R62 VSS.n22 VSS.n17 57.864
R63 VSS.n21 VSS.n20 15.3475
R64 VSS.n51 VSS.t24 12.5437
R65 VSS.n37 VSS.t3 12.4687
R66 VSS.n31 VSS.t22 12.4687
R67 VSS.n19 VSS.t18 12.4687
R68 VSS.n26 VSS.t5 12.4687
R69 VSS.n41 VSS.t16 12.4687
R70 VSS.n4 VSS.t10 12.4687
R71 VSS.n1 VSS.t13 12.4687
R72 VSS.n38 VSS.t8 12.4687
R73 VSS.n14 VSS.t20 12.4675
R74 VSS.n29 VSS.n28 11.6695
R75 VSS.n15 VSS.n14 10.4017
R76 VSS.n19 VSS.n18 10.4005
R77 VSS.n26 VSS.n25 10.4005
R78 VSS.n5 VSS.n4 10.4005
R79 VSS.n33 VSS.n1 10.4005
R80 VSS.n51 VSS.n50 10.4005
R81 VSS.n42 VSS.n41 10.4005
R82 VSS.n32 VSS.n31 10.4005
R83 VSS.n37 VSS.n36 10.4005
R84 VSS.n31 VSS.n0 9.86036
R85 VSS.n28 VSS.n27 6.42418
R86 VSS.n20 VSS.n19 6.02652
R87 VSS.n39 VSS.n38 5.75457
R88 VSS.n39 VSS.n2 5.48837
R89 VSS.n41 VSS.n40 5.44665
R90 VSS.n40 VSS.n37 5.3877
R91 VSS.n27 VSS.n26 4.66984
R92 VSS.n14 VSS.n12 4.6547
R93 VSS.n20 VSS.n12 1.34731
R94 VSS.n40 VSS.n39 1.2245
R95 VSS.n27 VSS.n12 1.03428
R96 VSS.n52 VSS.n2 0.820259
R97 VSS VSS.n0 0.783577
R98 VSS.n28 VSS.n0 0.664346
R99 VSS.n53 VSS.n52 0.652808
R100 VSS VSS.n53 0.348192
R101 VSS.n4 VSS.n2 0.323682
R102 VSS.n53 VSS.n1 0.322765
R103 VSS.n52 VSS.n51 0.314599
R104 a_n359_n5759.t8 a_n359_n5759.t5 69.3505
R105 a_n359_n5759.t4 a_n359_n5759.t3 69.3505
R106 a_n359_n5759.t6 a_n359_n5759.t7 53.4469
R107 a_n359_n5759.n2 a_n359_n5759.t6 35.2609
R108 a_n359_n5759.n1 a_n359_n5759.t8 30.3133
R109 a_n359_n5759.n2 a_n359_n5759.t4 25.048
R110 a_n359_n5759.t0 a_n359_n5759.n3 12.3005
R111 a_n359_n5759.n1 a_n359_n5759.n0 5.78668
R112 a_n359_n5759.n0 a_n359_n5759.t2 4.33383
R113 a_n359_n5759.n0 a_n359_n5759.t1 4.33383
R114 a_n359_n5759.n3 a_n359_n5759.n2 0.519935
R115 a_n359_n5759.n3 a_n359_n5759.n1 0.494983
R116 Q Q.t0 12.6202
R117 Q Q.t1 12.341
R118 VDD.n8 VDD.t23 715.11
R119 VDD.n11 VDD.t20 714.49
R120 VDD.n18 VDD.t21 713.694
R121 VDD.n14 VDD.t6 713.688
R122 VDD.n17 VDD.t18 713.688
R123 VDD.n12 VDD.t26 713.688
R124 VDD.n16 VDD.t8 713.688
R125 VDD.n9 VDD.t0 713.688
R126 VDD.n6 VDD.t4 713.688
R127 VDD.n0 VDD.t14 713.688
R128 VDD.n3 VDD.t2 713.688
R129 VDD.n2 VDD.t11 713.688
R130 VDD.t26 VDD.t16 434.784
R131 VDD.t0 VDD.t13 434.784
R132 VDD.t14 VDD.t24 434.784
R133 VDD.t2 VDD.t10 434.784
R134 VDD.n0 VDD.t25 13.7623
R135 VDD.n13 VDD.t17 12.5331
R136 VDD.n17 VDD.t19 12.1992
R137 VDD.n16 VDD.t9 12.1992
R138 VDD.n6 VDD.t5 12.1992
R139 VDD.n3 VDD.t3 12.1992
R140 VDD.n2 VDD.t12 12.1992
R141 VDD.n14 VDD.t7 12.198
R142 VDD.n10 VDD.t1 12.1968
R143 VDD.n18 VDD.t22 12.192
R144 VDD.n12 VDD.t27 12.1422
R145 VDD.n1 VDD.t15 12.1411
R146 VDD.n19 VDD.n18 11.4596
R147 VDD.n16 VDD.n15 9.90617
R148 VDD.n4 VDD.n2 7.0573
R149 VDD.n7 VDD.n5 5.46986
R150 VDD.n5 VDD.n1 5.05424
R151 VDD.n4 VDD.n3 5.0066
R152 VDD.n20 VDD.n19 3.429
R153 VDD.n11 VDD.n10 1.6793
R154 VDD.n19 VDD.n17 1.5236
R155 VDD.n9 VDD.n8 1.27962
R156 VDD.n13 VDD.n12 1.1387
R157 VDD VDD.n11 0.864995
R158 VDD.n5 VDD.n4 0.845079
R159 VDD.n20 VDD.n16 0.527474
R160 VDD.n15 VDD.n14 0.516611
R161 VDD.n15 VDD.n13 0.457423
R162 VDD.n8 VDD.n7 0.351026
R163 VDD VDD.n20 0.00545413
R164 VDD.n10 VDD.n9 0.00286842
R165 VDD.n7 VDD.n6 0.00168421
R166 VDD.n1 VDD.n0 0.00153448
R167 RSTN.t0 RSTN.t3 89.2951
R168 RSTN.t2 RSTN.t1 89.2951
R169 RSTN.n0 RSTN.t2 44.9198
R170 RSTN.n0 RSTN.t0 24.9469
R171 RSTN RSTN.n0 0.00286842
R172 D.t1 D.t0 53.4469
R173 D D.t1 24.9505
R174 CLK.t1 CLK.t0 69.3505
R175 CLK CLK.t1 24.9517
R176 Qb Qb.t0 12.6395
R177 Qb Qb.t1 12.3217
C0 VDD a_n1342_n5730# 1.71536f
C1 a_n249_n4912# a_881_n5758# 0.19693f
C2 a_n1374_n6642# a_n1342_n5730# 1.67868f
C3 RSTN a_n249_n4912# 0.28644f
C4 a_n249_n4912# a_n1342_n5730# 0.21283f
C5 a_1056_n4015# a_881_n5758# 0.25267f
C6 VDD a_991_n4911# 0.76938f
C7 a_881_n5758# a_n1342_n5730# 0.31376f
C8 a_n1374_n6642# a_991_n4911# 0.22275f
C9 VDD D 0.18707f
C10 VDD a_n912_n3722# 0.83176f
C11 a_n249_n4912# a_991_n4911# 0.11019f
C12 VDD CLK 0.28794f
C13 VDD a_n1374_n6642# 1.886f
C14 VDD a_n249_n4912# 0.56511f
C15 a_991_n4911# a_881_n5758# 0.35092f
C16 a_n1374_n6642# a_n249_n4912# 0.23084f
C17 a_1056_n4015# a_991_n4911# 0.10365f
C18 VDD a_881_n5758# 1.18904f
C19 RSTN a_991_n4911# 0.29193f
C20 VDD a_1056_n4015# 0.95856f
C21 a_n1374_n6642# a_881_n5758# 0.24946f
C22 VDD Qb 0.10704f
C23 VDD RSTN 0.80322f
C24 a_n1374_n6642# a_1056_n4015# 0.2678f
C25 Q VSS 0.25589f
C26 CLK VSS 0.39888f
C27 RSTN VSS 1.32962f
C28 D VSS 0.27844f
C29 Qb VSS 0.15428f
C30 VDD VSS 18.83505f
C31 a_991_n4911# VSS 1.33038f
C32 a_n249_n4912# VSS 2.53842f
C33 a_881_n5758# VSS 0.89126f
C34 a_1056_n4015# VSS 1.26966f
C35 a_n1374_n6642# VSS 5.44569f
C36 a_n1342_n5730# VSS 6.88765f
C37 a_n912_n3722# VSS 0.62392f
C38 VDD.n8 VSS 0.11133f
C39 VDD.n11 VSS 0.13113f
C40 VDD.n19 VSS 0.21025f
C41 VDD.n20 VSS 0.10843f
C42 a_n359_n5759.t8 VSS 0.19196f
C43 a_n359_n5759.n1 VSS 1.35777f
C44 a_n359_n5759.t6 VSS 0.11284f
C45 a_n359_n5759.n2 VSS 0.45569f
C46 a_n359_n5759.n3 VSS 0.14466f
.ends

