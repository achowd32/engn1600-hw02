* Extracted by KLayout with GF180MCU LVS runset on : 14/02/2026 05:24

.SUBCKT TGATE vss VDD IN OUT C CBAR
M$1 OUT CBAR IN VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$2 OUT C IN vss nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U PD=2.1U
.ENDS TGATE
