* Extracted by KLayout with GF180MCU LVS runset on : 22/02/2026 22:49

.SUBCKT dff VSS Q CLK VDD RSTN Qb D
M$1 VDD \$1 \$17 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$2 VDD \$7 Q VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$3 \$19 \$7 \$5 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$4 \$19 \$17 VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$5 \$5 \$1 \$9 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$6 VDD CLK \$1 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$7 \$7 \$5 VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$8 \$7 RSTN VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$9 \$22 \$9 VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$10 \$22 RSTN VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$11 VDD \$34 \$9 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$12 \$22 \$1 \$34 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$13 \$49 D \$34 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$14 \$49 \$17 VDD VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.1092P PS=2.18U
+ PD=0.94U
M$15 VDD \$7 \$42 VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$16 VDD \$42 Qb VDD pfet_03v3 L=0.28U W=0.42U AS=0.2822P AD=0.2822P PS=2.18U
+ PD=2.18U
M$17 VSS \$1 \$17 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2625P AD=0.2667P PS=2.09U
+ PD=2.11U
M$18 VSS \$7 Q VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$19 \$12 \$7 \$5 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$20 \$12 \$1 VSS VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$21 \$5 \$17 \$9 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$22 VSS CLK \$1 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$23 \$27 \$5 \$7 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$24 \$27 RSTN VSS VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$25 \$28 \$9 \$22 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$26 \$28 RSTN VSS VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$27 VSS \$34 \$9 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$28 \$22 \$17 \$34 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$29 \$47 D \$34 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$30 \$47 \$1 VSS VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.1092P PS=2.1U
+ PD=0.94U
M$31 VSS \$7 \$42 VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
M$32 VSS \$42 Qb VSS nfet_03v3 L=0.28U W=0.42U AS=0.2646P AD=0.2646P PS=2.1U
+ PD=2.1U
.ENDS dff
