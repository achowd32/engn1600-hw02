** sch_path: /foss/designs/CAD2/nand2.sch
.subckt nand2 vdd OUT IN0 IN1 vss
*.PININFO IN0:I IN1:I OUT:O vdd:B vss:B
M1 net1 IN1 vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M3 OUT IN0 vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M4 OUT IN1 vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M2 OUT IN0 net1 vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
.ends
