* NGSPICE file created from dff_flat.ext - technology: gf180mcuD

.subckt dff_flat CHECK VDD CLK RSTN VSS D Q Qb
X0 a_n249_n4912# a_n1374_n6642# RSTN.t2 VSS.t12 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X1 VSS.t4 a_n359_n5759.t3 Q.t1 VSS.t3 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X2 a_n359_n5759.t1 a_n249_n4912# VDD.t23 VDD.t22 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X3 VDD.t8 a_n89_n4912# a_881_n5758# VDD.t7 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X4 VDD.t17 a_n1374_n6642# a_1067_n6116# VDD.t16 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X5 a_2281_n4424# D.t0 CHECK.t3 VSS.t19 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X6 VSS.t6 CLK.t0 a_n1342_n5730# VSS.t5 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X7 a_2280_n3998# D.t1 CHECK.t2 VDD.t4 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X8 VDD.t1 CLK.t1 a_n1342_n5730# VDD.t0 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X9 VSS.t18 a_n1342_n5730# a_n1374_n6642# VSS.t17 nfet_03v3 ad=0.2667p pd=2.11u as=0.2625p ps=2.09u w=0.42u l=0.28u
X10 a_1059_n5756# RSTN.t4 a_881_n5758# VSS.t23 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X11 VSS.t1 CHECK.t4 RSTN.t0 VSS.t0 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X12 VSS.t16 a_n1342_n5730# a_1068_n6542# VSS.t15 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X13 VSS.t25 a_n912_n3722# Qb.t1 VSS.t24 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X14 VSS.t10 a_n89_n4912# a_n181_n5757# VSS.t9 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X15 VDD.t13 a_n359_n5759.t4 Q.t0 VDD.t12 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X16 a_n249_n4912# a_n1342_n5730# RSTN.t3 VDD.t21 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X17 VSS.t22 a_n359_n5759.t5 a_n912_n3722# VSS.t21 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X18 VDD.t20 a_n1342_n5730# a_n1374_n6642# VDD.t19 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X19 a_881_n5758# a_n1374_n6642# CHECK.t0 VSS.t11 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
X20 VDD.t27 a_n912_n3722# Qb.t0 VDD.t26 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X21 VSS.t14 a_n1342_n5730# a_2281_n4424# VSS.t13 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X22 VDD.t6 a_n89_n4912# a_n359_n5759.t0 VDD.t5 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X23 VDD.t15 a_n1374_n6642# a_2280_n3998# VDD.t14 pfet_03v3 ad=0.2822p pd=2.18u as=0.1092p ps=0.94u w=0.42u l=0.28u
X24 a_1067_n6116# a_n359_n5759.t6 a_n249_n4912# VDD.t11 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X25 a_881_n5758# RSTN.t5 VDD.t25 VDD.t24 pfet_03v3 ad=0.1092p pd=0.94u as=0.2822p ps=2.18u w=0.42u l=0.28u
X26 VSS.t8 a_n89_n4912# a_1059_n5756# VSS.t7 nfet_03v3 ad=0.2646p pd=2.1u as=0.1092p ps=0.94u w=0.42u l=0.28u
X27 VDD.t3 CHECK.t5 RSTN.t1 VDD.t2 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X28 a_881_n5758# a_n1342_n5730# CHECK.t1 VDD.t18 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
X29 a_1068_n6542# a_n359_n5759.t7 a_n249_n4912# VSS.t2 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X30 a_n181_n5757# a_n249_n4912# a_n359_n5759.t2 VSS.t20 nfet_03v3 ad=0.1092p pd=0.94u as=0.2646p ps=2.1u w=0.42u l=0.28u
X31 VDD.t10 a_n359_n5759.t8 a_n912_n3722# VDD.t9 pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
R0 RSTN.t5 RSTN.n3 72.3487
R1 RSTN RSTN.t5 24.9493
R2 RSTN.n3 RSTN.t4 16.9469
R3 RSTN.n1 RSTN.t2 12.9962
R4 RSTN.n0 RSTN.t1 12.66
R5 RSTN.n0 RSTN.t0 12.3135
R6 RSTN.n1 RSTN.t3 12.0263
R7 RSTN.n3 RSTN.n2 9.90023
R8 RSTN.n2 RSTN.n1 0.39464
R9 RSTN.n2 RSTN.n0 0.156576
R10 VSS.n23 VSS.n16 749278
R11 VSS.n16 VSS.t19 91327.6
R12 VSS.n5 VSS.n3 64653.5
R13 VSS.n50 VSS.n3 47027.8
R14 VSS.n13 VSS.n8 11150.5
R15 VSS.t24 VSS.n46 10656.3
R16 VSS.n46 VSS.n45 9310.54
R17 VSS.n6 VSS.n3 9172.39
R18 VSS.n17 VSS.n8 8859.18
R19 VSS.n46 VSS.n7 7710.44
R20 VSS.n43 VSS.n9 6769.51
R21 VSS.n35 VSS.n34 6625.47
R22 VSS.n45 VSS.n8 5874.35
R23 VSS.t17 VSS.n49 4464.13
R24 VSS.n13 VSS.n11 4354.26
R25 VSS.n30 VSS.n10 4226.8
R26 VSS.n29 VSS.n11 4102.23
R27 VSS.n45 VSS.n44 3676.98
R28 VSS.n24 VSS.n23 3564.92
R29 VSS.n44 VSS.t11 2894.81
R30 VSS.n47 VSS.n7 2588.74
R31 VSS.t3 VSS.n3 2474.65
R32 VSS.n49 VSS.n48 2224.45
R33 VSS.n49 VSS.t5 1774.36
R34 VSS.n48 VSS.n6 1755.92
R35 VSS.n22 VSS.n21 1702.15
R36 VSS.t0 VSS.n24 1689.9
R37 VSS.n24 VSS.n10 1589.78
R38 VSS.t5 VSS.n5 1493.57
R39 VSS.t13 VSS.n15 1430.46
R40 VSS.n25 VSS.t0 1413.04
R41 VSS.t23 VSS.n9 1360.03
R42 VSS.n21 VSS.t11 1205.49
R43 VSS.t21 VSS.n7 1196.19
R44 VSS.n48 VSS.n47 1177.13
R45 VSS.n18 VSS.t7 1172.44
R46 VSS.n23 VSS.n22 1095.11
R47 VSS.n25 VSS.n11 1090.87
R48 VSS.n36 VSS.t9 1070.49
R49 VSS.n34 VSS.t2 1055.67
R50 VSS.n42 VSS.t21 992.063
R51 VSS.n30 VSS.t12 940.115
R52 VSS.n50 VSS.t17 920.712
R53 VSS.t19 VSS.t13 915.494
R54 VSS.n18 VSS.n10 900.433
R55 VSS.n34 VSS.n33 836.077
R56 VSS.n36 VSS.n35 822.135
R57 VSS.n32 VSS.n30 797.649
R58 VSS.t7 VSS.t23 750.361
R59 VSS.t9 VSS.t20 685.112
R60 VSS.n17 VSS.n16 674.74
R61 VSS.n38 VSS.n7 671.655
R62 VSS.n43 VSS.n42 615.08
R63 VSS.n33 VSS.t3 604.99
R64 VSS.t15 VSS.n32 576.241
R65 VSS.t12 VSS.n29 492.724
R66 VSS.n44 VSS.n43 472.2
R67 VSS.n15 VSS.n13 469.19
R68 VSS.t20 VSS.n6 466.733
R69 VSS.n47 VSS.t24 415.238
R70 VSS.t2 VSS.t15 368.795
R71 VSS.n35 VSS.n9 317.529
R72 VSS.n22 VSS.n17 57.864
R73 VSS.n21 VSS.n20 15.3475
R74 VSS.n51 VSS.t18 12.5437
R75 VSS.n37 VSS.t10 12.4687
R76 VSS.n31 VSS.t16 12.4687
R77 VSS.n19 VSS.t8 12.4687
R78 VSS.n26 VSS.t1 12.4687
R79 VSS.n41 VSS.t22 12.4687
R80 VSS.n4 VSS.t6 12.4687
R81 VSS.n1 VSS.t4 12.4687
R82 VSS.n38 VSS.t25 12.4687
R83 VSS.n14 VSS.t14 12.4675
R84 VSS.n29 VSS.n28 11.6695
R85 VSS.n15 VSS.n14 10.4017
R86 VSS.n19 VSS.n18 10.4005
R87 VSS.n26 VSS.n25 10.4005
R88 VSS.n5 VSS.n4 10.4005
R89 VSS.n33 VSS.n1 10.4005
R90 VSS.n51 VSS.n50 10.4005
R91 VSS.n42 VSS.n41 10.4005
R92 VSS.n32 VSS.n31 10.4005
R93 VSS.n37 VSS.n36 10.4005
R94 VSS.n31 VSS.n0 9.86036
R95 VSS.n28 VSS.n27 6.42418
R96 VSS.n20 VSS.n19 6.02652
R97 VSS.n39 VSS.n38 5.75457
R98 VSS.n39 VSS.n2 5.48837
R99 VSS.n41 VSS.n40 5.44665
R100 VSS.n40 VSS.n37 5.3877
R101 VSS.n27 VSS.n26 4.66984
R102 VSS.n14 VSS.n12 4.6547
R103 VSS.n20 VSS.n12 1.34731
R104 VSS.n40 VSS.n39 1.2245
R105 VSS.n27 VSS.n12 1.03428
R106 VSS.n52 VSS.n2 0.820259
R107 VSS VSS.n0 0.783577
R108 VSS.n28 VSS.n0 0.664346
R109 VSS.n53 VSS.n52 0.652808
R110 VSS VSS.n53 0.348192
R111 VSS.n4 VSS.n2 0.323682
R112 VSS.n53 VSS.n1 0.322765
R113 VSS.n52 VSS.n51 0.314599
R114 a_n359_n5759.t8 a_n359_n5759.t5 69.3505
R115 a_n359_n5759.t4 a_n359_n5759.t3 69.3505
R116 a_n359_n5759.t6 a_n359_n5759.t7 53.4469
R117 a_n359_n5759.n0 a_n359_n5759.t6 35.2609
R118 a_n359_n5759.n2 a_n359_n5759.t8 30.3133
R119 a_n359_n5759.n0 a_n359_n5759.t4 25.048
R120 a_n359_n5759.n1 a_n359_n5759.t2 12.3005
R121 a_n359_n5759.n3 a_n359_n5759.n2 5.78668
R122 a_n359_n5759.t0 a_n359_n5759.n3 4.33383
R123 a_n359_n5759.n3 a_n359_n5759.t1 4.33383
R124 a_n359_n5759.n1 a_n359_n5759.n0 0.519935
R125 a_n359_n5759.n2 a_n359_n5759.n1 0.494983
R126 Q Q.t1 12.6202
R127 Q Q.t0 12.341
R128 VDD.n8 VDD.t21 715.11
R129 VDD.n11 VDD.t18 714.49
R130 VDD.n18 VDD.t19 713.694
R131 VDD.n14 VDD.t26 713.688
R132 VDD.n17 VDD.t0 713.688
R133 VDD.n12 VDD.t5 713.688
R134 VDD.n16 VDD.t9 713.688
R135 VDD.n9 VDD.t14 713.688
R136 VDD.n6 VDD.t2 713.688
R137 VDD.n0 VDD.t7 713.688
R138 VDD.n3 VDD.t16 713.688
R139 VDD.n2 VDD.t12 713.688
R140 VDD.t5 VDD.t22 434.784
R141 VDD.t14 VDD.t4 434.784
R142 VDD.t7 VDD.t24 434.784
R143 VDD.t16 VDD.t11 434.784
R144 VDD.n0 VDD.t25 13.7623
R145 VDD.n13 VDD.t23 12.5331
R146 VDD.n17 VDD.t1 12.1992
R147 VDD.n16 VDD.t10 12.1992
R148 VDD.n6 VDD.t3 12.1992
R149 VDD.n3 VDD.t17 12.1992
R150 VDD.n2 VDD.t13 12.1992
R151 VDD.n14 VDD.t27 12.198
R152 VDD.n10 VDD.t15 12.1968
R153 VDD.n18 VDD.t20 12.192
R154 VDD.n12 VDD.t6 12.1422
R155 VDD.n1 VDD.t8 12.1411
R156 VDD.n19 VDD.n18 11.4596
R157 VDD.n16 VDD.n15 9.90617
R158 VDD.n4 VDD.n2 7.0573
R159 VDD.n7 VDD.n5 5.46986
R160 VDD.n5 VDD.n1 5.05424
R161 VDD.n4 VDD.n3 5.0066
R162 VDD.n20 VDD.n19 3.429
R163 VDD.n11 VDD.n10 1.6793
R164 VDD.n19 VDD.n17 1.5236
R165 VDD.n9 VDD.n8 1.27962
R166 VDD.n13 VDD.n12 1.1387
R167 VDD VDD.n11 0.864995
R168 VDD.n5 VDD.n4 0.845079
R169 VDD.n20 VDD.n16 0.527474
R170 VDD.n15 VDD.n14 0.516611
R171 VDD.n15 VDD.n13 0.457423
R172 VDD.n8 VDD.n7 0.351026
R173 VDD VDD.n20 0.00545413
R174 VDD.n10 VDD.n9 0.00286842
R175 VDD.n7 VDD.n6 0.00168421
R176 VDD.n1 VDD.n0 0.00153448
R177 D.t1 D.t0 53.4469
R178 D D.t1 24.9505
R179 CHECK.t5 CHECK.t4 69.3505
R180 CHECK.n1 CHECK.t5 25.414
R181 CHECK.n0 CHECK.t1 12.667
R182 CHECK CHECK.t2 12.3758
R183 CHECK.n2 CHECK.t3 12.3005
R184 CHECK.n0 CHECK.t0 12.3005
R185 CHECK.n1 CHECK.n0 1.9362
R186 CHECK.n2 CHECK.n1 0.19099
R187 CHECK CHECK.n2 0.179078
R188 CLK.t1 CLK.t0 69.3505
R189 CLK CLK.t1 24.9517
R190 Qb Qb.t1 12.6395
R191 Qb Qb.t0 12.3217
C0 RSTN CHECK 0.10365f
C1 VDD a_n89_n4912# 0.80322f
C2 a_n1342_n5730# a_881_n5758# 0.31376f
C3 a_n249_n4912# VDD 0.56511f
C4 a_n1374_n6642# a_n249_n4912# 0.23084f
C5 RSTN VDD 0.76938f
C6 a_n249_n4912# a_n89_n4912# 0.28644f
C7 a_881_n5758# CHECK 0.25267f
C8 RSTN a_n1374_n6642# 0.22275f
C9 RSTN a_n89_n4912# 0.29193f
C10 VDD a_n1342_n5730# 1.71536f
C11 RSTN a_n249_n4912# 0.11019f
C12 a_n1374_n6642# a_n1342_n5730# 1.67868f
C13 VDD a_881_n5758# 1.18904f
C14 CLK VDD 0.28794f
C15 a_n1374_n6642# a_881_n5758# 0.24946f
C16 VDD CHECK 0.95856f
C17 a_n249_n4912# a_n1342_n5730# 0.21283f
C18 a_n1374_n6642# CHECK 0.2678f
C19 a_n912_n3722# VDD 0.83176f
C20 a_n249_n4912# a_881_n5758# 0.19693f
C21 Qb VDD 0.10704f
C22 RSTN a_881_n5758# 0.35092f
C23 a_n1374_n6642# VDD 1.886f
C24 VDD D 0.18707f
C25 Q VSS 0.25589f
C26 CLK VSS 0.39888f
C27 RSTN VSS 1.33038f
C28 CHECK VSS 1.26966f
C29 D VSS 0.27844f
C30 Qb VSS 0.15428f
C31 VDD VSS 18.83505f
C32 a_n89_n4912# VSS 1.32962f
C33 a_n249_n4912# VSS 2.53842f
C34 a_881_n5758# VSS 0.89126f
C35 a_n1374_n6642# VSS 5.44569f
C36 a_n1342_n5730# VSS 6.88765f
C37 a_n912_n3722# VSS 0.62392f
C38 VDD.n8 VSS 0.11133f
C39 VDD.n11 VSS 0.13113f
C40 VDD.n19 VSS 0.21025f
C41 VDD.n20 VSS 0.10843f
C42 a_n359_n5759.t8 VSS 0.19196f
C43 a_n359_n5759.t6 VSS 0.11284f
C44 a_n359_n5759.n0 VSS 0.45569f
C45 a_n359_n5759.n1 VSS 0.14466f
C46 a_n359_n5759.n2 VSS 1.35777f
.ends

